* NGSPICE file created from pes_decoder.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

.subckt pes_decoder VGND VPWR clk in[0] in[1] in[2] out[0] out[1] out[2] out[3] out[4]
+ out[5] out[6] out[7]
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput7 net7 VGND VGND VPWR VPWR out[3] sky130_fd_sc_hd__buf_1
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xout_sky130_fd_sc_hd__nor4b_2_Y net1 net2 net3 clknet_1_1__leaf_clk VGND VGND VPWR
+ VPWR net4 sky130_fd_sc_hd__nor4b_2
XFILLER_0_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput10 net10 VGND VGND VPWR VPWR out[6] sky130_fd_sc_hd__buf_1
Xoutput8 net8 VGND VGND VPWR VPWR out[4] sky130_fd_sc_hd__buf_1
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR out[5] sky130_fd_sc_hd__buf_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput11 net11 VGND VGND VPWR VPWR out[7] sky130_fd_sc_hd__buf_1
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclk_sky130_fd_sc_hd__and4_2_D net1 net2 net3 clknet_1_1__leaf_clk VGND VGND VPWR
+ VPWR out_sky130_fd_sc_hd__buf_1_X_A sky130_fd_sc_hd__and4_2
XFILLER_0_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclk_sky130_fd_sc_hd__and4b_2_B net3 clknet_1_1__leaf_clk net1 net2 VGND VGND VPWR
+ VPWR clk_sky130_fd_sc_hd__and4b_2_B_X sky130_fd_sc_hd__and4b_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclk_sky130_fd_sc_hd__and4b_2_C net2 net3 clknet_1_0__leaf_clk net1 VGND VGND VPWR
+ VPWR clk_sky130_fd_sc_hd__and4b_2_C_X sky130_fd_sc_hd__and4b_2
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclk_sky130_fd_sc_hd__and4b_2_D net1 net2 net3 clknet_1_0__leaf_clk VGND VGND VPWR
+ VPWR clk_sky130_fd_sc_hd__and4b_2_D_X sky130_fd_sc_hd__and4b_2
XFILLER_0_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 in[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 in[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclk_sky130_fd_sc_hd__and4bb_2_C net1 net3 clknet_1_1__leaf_clk net2 VGND VGND VPWR
+ VPWR out_sky130_fd_sc_hd__buf_1_X_5_A sky130_fd_sc_hd__and4bb_2
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclk_sky130_fd_sc_hd__and4bb_2_D net1 net2 net3 clknet_1_0__leaf_clk VGND VGND VPWR
+ VPWR out_sky130_fd_sc_hd__buf_1_X_3_A sky130_fd_sc_hd__and4bb_2
XFILLER_0_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xout_sky130_fd_sc_hd__buf_1_X out_sky130_fd_sc_hd__buf_1_X_A VGND VGND VPWR VPWR net11
+ sky130_fd_sc_hd__buf_1
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xout_sky130_fd_sc_hd__buf_1_X_1 clk_sky130_fd_sc_hd__and4b_2_D_X VGND VGND VPWR VPWR
+ net10 sky130_fd_sc_hd__buf_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xout_sky130_fd_sc_hd__buf_1_X_2 clk_sky130_fd_sc_hd__and4b_2_C_X VGND VGND VPWR VPWR
+ net9 sky130_fd_sc_hd__buf_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xout_sky130_fd_sc_hd__buf_1_X_3 out_sky130_fd_sc_hd__buf_1_X_3_A VGND VGND VPWR VPWR
+ net8 sky130_fd_sc_hd__buf_1
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclk_sky130_fd_sc_hd__and4bb_2_C_1 net2 net3 clknet_1_0__leaf_clk net1 VGND VGND VPWR
+ VPWR out_sky130_fd_sc_hd__buf_1_X_6_A sky130_fd_sc_hd__and4bb_2
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xout_sky130_fd_sc_hd__buf_1_X_4 clk_sky130_fd_sc_hd__and4b_2_B_X VGND VGND VPWR VPWR
+ net7 sky130_fd_sc_hd__buf_1
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xout_sky130_fd_sc_hd__buf_1_X_5 out_sky130_fd_sc_hd__buf_1_X_5_A VGND VGND VPWR VPWR
+ net6 sky130_fd_sc_hd__buf_1
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xout_sky130_fd_sc_hd__buf_1_X_6 out_sky130_fd_sc_hd__buf_1_X_6_A VGND VGND VPWR VPWR
+ net5 sky130_fd_sc_hd__buf_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR out[0] sky130_fd_sc_hd__buf_1
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR out[1] sky130_fd_sc_hd__buf_1
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput6 net6 VGND VGND VPWR VPWR out[2] sky130_fd_sc_hd__buf_1
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

