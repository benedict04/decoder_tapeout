magic
tech sky130A
magscale 1 2
timestamp 1700889145
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37584
<< metal2 >>
rect 662 39200 718 40000
rect 13542 39200 13598 40000
rect 26422 39200 26478 40000
rect 39302 39200 39358 40000
rect 18 0 74 800
rect 12898 0 12954 800
rect 25778 0 25834 800
rect 38658 0 38714 800
<< obsm2 >>
rect 20 39144 606 39200
rect 774 39144 13486 39200
rect 13654 39144 26366 39200
rect 26534 39144 39246 39200
rect 20 856 39356 39144
rect 130 800 12842 856
rect 13010 800 25722 856
rect 25890 800 38602 856
rect 38770 800 39356 856
<< metal3 >>
rect 0 27208 800 27328
rect 39200 25848 40000 25968
rect 0 13608 800 13728
rect 39200 12248 40000 12368
<< obsm3 >>
rect 800 27408 39200 37569
rect 880 27128 39200 27408
rect 800 26048 39200 27128
rect 800 25768 39120 26048
rect 800 13808 39200 25768
rect 880 13528 39200 13808
rect 800 12448 39200 13528
rect 800 12168 39120 12448
rect 800 2143 39200 12168
<< metal4 >>
rect 1944 2128 2264 37584
rect 2604 2128 2924 37584
rect 6944 2128 7264 37584
rect 7604 2128 7924 37584
rect 11944 2128 12264 37584
rect 12604 2128 12924 37584
rect 16944 2128 17264 37584
rect 17604 2128 17924 37584
rect 21944 2128 22264 37584
rect 22604 2128 22924 37584
rect 26944 2128 27264 37584
rect 27604 2128 27924 37584
rect 31944 2128 32264 37584
rect 32604 2128 32924 37584
rect 36944 2128 37264 37584
rect 37604 2128 37924 37584
<< metal5 >>
rect 1056 33676 38872 33996
rect 1056 33016 38872 33336
rect 1056 28676 38872 28996
rect 1056 28016 38872 28336
rect 1056 23676 38872 23996
rect 1056 23016 38872 23336
rect 1056 18676 38872 18996
rect 1056 18016 38872 18336
rect 1056 13676 38872 13996
rect 1056 13016 38872 13336
rect 1056 8676 38872 8996
rect 1056 8016 38872 8336
rect 1056 3676 38872 3996
rect 1056 3016 38872 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 38872 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 38872 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 38872 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18676 38872 18996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 23676 38872 23996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 28676 38872 28996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 33676 38872 33996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 38872 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 38872 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 38872 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18016 38872 18336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23016 38872 23336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 28016 38872 28336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 33016 38872 33336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 13608 800 13728 6 clk
port 3 nsew signal input
rlabel metal2 s 39302 39200 39358 40000 6 in[0]
port 4 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 in[1]
port 5 nsew signal input
rlabel metal2 s 18 0 74 800 6 in[2]
port 6 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 out[0]
port 7 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 out[1]
port 8 nsew signal output
rlabel metal2 s 26422 39200 26478 40000 6 out[2]
port 9 nsew signal output
rlabel metal3 s 39200 25848 40000 25968 6 out[3]
port 10 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 out[4]
port 11 nsew signal output
rlabel metal2 s 662 39200 718 40000 6 out[5]
port 12 nsew signal output
rlabel metal2 s 13542 39200 13598 40000 6 out[6]
port 13 nsew signal output
rlabel metal3 s 39200 12248 40000 12368 6 out[7]
port 14 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 927580
string GDS_FILE /home/hardhik/decoder_tapeout/openlane/pes_decoder/runs/23_11_25_00_11/results/signoff/pes_decoder.magic.gds
string GDS_START 75164
<< end >>

